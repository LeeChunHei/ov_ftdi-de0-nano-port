module test_ft245_sync(
	input		CLOCK_50,
	output	[7:0]LED,
	output	[2:0]leds,
	input		ftdi_clk,
	output	[7:0]ftdi_d__,
	output	ftdi_rxf_n__,
	output	ftdi_txe_n__,
	output	ftdi_rd_n__,
	output	ftdi_wr_n__,
	output	ftdi_siwua_n__,
	output	ftdi_oe_n__,
	output	fifo_rinc__,
	output	[7:0]fifo_rdata__,
	output	fifo_rempty__,
	output	fifo_winc__,
	output	[7:0]fifo_wdata__,
	output	fifo_wfull__,
	output	fifo_tx_ind__,
	output	fifo_rx_ind__
);

	wire pll_rst;
	wire pll_locked;
	wire sys_clk;
	wire sys_rst_n;
	
	
	wire	[7:0]ftdi_d;
	reg	[7:0]ftdi_d_reg;
	reg	ftdi_d_oe;
	reg	_ftdi_rxf_n;
	reg	_ftdi_txe_n;
	wire	ftdi_rd_n;
	wire	ftdi_wr_n;
	wire	ftdi_siwua_n;
	wire	ftdi_oe_n;
	reg	fifo_rinc;
	wire	[7:0]fifo_rdata;
	wire	fifo_rempty;
	reg	fifo_winc;
	reg	[7:0]fifo_wdata;
	wire	fifo_wfull;
	wire	fifo_tx_ind;
	wire	fifo_rx_ind;
	
	assign pll_rst = 0;
	assign sys_rst_n = pll_locked;
	
	assign ftdi_d = ftdi_d_oe ? ftdi_d_reg : 8'bzzzzzzzz;
	assign ftdi_d__ = ftdi_d;
	assign ftdi_rxf_n__ = _ftdi_rxf_n;
	assign ftdi_txe_n__ = _ftdi_txe_n;
	assign ftdi_rd_n__ = ftdi_rd_n;
	assign ftdi_wr_n__ = ftdi_wr_n;
	assign ftdi_siwua_n__ = ftdi_siwua_n;
	assign ftdi_oe_n__ = ftdi_oe_n;
	assign fifo_rinc__ = fifo_rinc;
	assign fifo_rdata__ = fifo_rdata;
	assign fifo_rempty__ = fifo_rempty;
	assign fifo_winc__ = fifo_winc;
	assign fifo_wdata__ = fifo_wdata;
	assign fifo_wfull__ = fifo_wfull;
	assign fifo_tx_ind__ = fifo_tx_ind;
	assign fifo_rx_ind__ = fifo_rx_ind;
	
	pll pll_0(
		.areset(pll_rst),
		.inclk0(CLOCK_50),
		.c0(sys_clk),
		.locked(pll_locked));
	
	syncFT245 ft245_bus(
		.io_clk(ftdi_clk),
		.io_d(ftdi_d),
		.io_rxf_n(_ftdi_rxf_n),
		.io_txe_n(_ftdi_txe_n),
		.io_rd_n(ftdi_rd_n),
		.io_wr_n(ftdi_wr_n),
		.io_siwua_n(ftdi_siwua_n),
		.io_oe_n(ftdi_oe_n),
		.rst_n(sys_rst_n),
		.sys_clk(sys_clk),
		.rinc(fifo_rinc),
		.rdata(fifo_rdata),
		.rempty(fifo_rempty),
		.winc(fifo_winc),
		.wdata(fifo_wdata),
		.wfull(fifo_wfull),
		.tx_ind(fifo_tx_ind),
		.rx_ind(fifo_rx_ind)
	);
	
	reg [7:0]ft_state;
	reg [7:0]ft_next_state;
	reg [7:0]count;
	
	reg [7:0]state;
	reg [7:0]next_state;
	
	parameter IDLE = 0;
	parameter WRITE0 = 1;
	parameter WRITE1 = 2;
	parameter WRITE2 = 3;
	parameter WRITE3 = 4;
	parameter WRITE4 = 5;
	parameter READ0 = 6;
	parameter READ1 = 7;
	parameter READ2 = 8;
	parameter READ3 = 9;
	parameter READ4 = 10;	
	
	always @(posedge ftdi_clk or negedge sys_rst_n) begin
		if (!sys_rst_n) begin
			ftdi_d_oe <= 0;
			_ftdi_rxf_n <= 1;
			_ftdi_txe_n <= 1;
			count <= 1;
			ft_state <= IDLE;
			ft_next_state <= IDLE;
		end
		else begin
			ft_state <= ft_next_state;
			case (ft_state)
				IDLE: begin
					ftdi_d_oe <= 0;
					_ftdi_rxf_n <= 1;
					_ftdi_txe_n <= 1;
					ft_next_state <= WRITE0;
				end
				WRITE0: begin
					_ftdi_rxf_n <= 0;
					ft_next_state <= WRITE1;
				end
				WRITE1: begin
					if (!ftdi_oe_n) begin
						count <= count + 1;
						ftdi_d_reg <= count;
						ftdi_d_oe <= 1;
						ft_next_state <= WRITE2;
					end
				end
				WRITE2: begin
					if (!ftdi_rd_n) begin
						count <= count + 1;
						ftdi_d_reg <= count;
						ftdi_d_oe <= 1;
					end
					if (ftdi_oe_n) begin
						ft_next_state <= WRITE3;
					end
					if (count > 2) begin
						_ftdi_rxf_n <= 1;
					end
				end
				WRITE3: begin
					ftdi_d_oe <= 0;
					ft_next_state <= IDLE;
				end
			endcase
		end
	end
	
	always @(posedge sys_clk or negedge sys_rst_n) begin
		if (!sys_rst_n) begin
			fifo_rinc <= 0;
			fifo_winc <= 0;
			fifo_wdata <= 0;
			state <= IDLE;
			next_state <= IDLE;
		end
		else begin
			if (!fifo_rempty) begin
				fifo_rinc <= 1;
			end
			else begin
				fifo_rinc <= 0;
			end
		
			state <= next_state;
//			case (ft_state)
//				IDLE: begin
//					ftdi_rxf_n <= 1;
//					ftdi_txe_n <= 1;
//					fifo_rinc <= 0;
//					fifo_winc <= 0;
//					fifo_wdata <= 0;
//				end
//			endcase
		end
	end
	
endmodule